// this a line compent
//
//


/*
 *
 * why
 */

// 中文你认得吗？？

module  

iopad
    (
        output  wire    [DW-1:0]    din,
        input   reg [DW-1:0]    dout,
`ifdef aa
        input   tri [DW-1:0]    dout_en,
`endif
        input clk,
        input   rst_n,
    );

